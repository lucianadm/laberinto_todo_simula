library verilog;
use verilog.vl_types.all;
entity pru_vlg_vec_tst is
end pru_vlg_vec_tst;
