library verilog;
use verilog.vl_types.all;
entity matriz_pru_vlg_check_tst is
    port(
        C0              : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end matriz_pru_vlg_check_tst;
