library verilog;
use verilog.vl_types.all;
entity actualiza_actual_vlg_vec_tst is
end actualiza_actual_vlg_vec_tst;
