library verilog;
use verilog.vl_types.all;
entity casillero_vlg_vec_tst is
end casillero_vlg_vec_tst;
