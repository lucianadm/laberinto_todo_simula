library verilog;
use verilog.vl_types.all;
entity matriz_pru_vlg_vec_tst is
end matriz_pru_vlg_vec_tst;
